
signature sMallocStatics {
	size_t getMaxSize(void);
	size_t getUsableSize(void);
	size_t getUsedSize(void);
	size_t getMallocSize(void);
	size_t getFreeSize(void);
	size_t getReallocSize(void);
};
