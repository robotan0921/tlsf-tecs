import( <sMalloc.cdl> );
import( "tTLSFStatics.cdl" );   //TODO: "" -> <>
import( <kernel.cdl> );

celltype tTLSFMalloc {
    // [inline]
        entry  sMalloc  eMalloc;
    entry   sMallocStatics  eMallocStatics;
    attr {
        /* memory pool size in bytes */
        size_t  memoryPoolSize;
    };
    var {
        [size_is( memoryPoolSize/ 8 )]
            uint64_t   *pool;
        size_t mallocSize;
        size_t freeSize;
        size_t reallocSize;
    };
};
