import( <sMalloc.cdl> );
import( <sMallocStatistics.cdl> );
import( <kernel.cdl> );

celltype tTLSFMalloc {
    [inline]
        entry  sMalloc  eMalloc;
    [inline]
        entry  sMallocStatistics    eMallocStatistics;
    attr {
        /* memory pool size in bytes */
        size_t  memoryPoolSize;
    };
    var {
        [size_is( memoryPoolSize/ 8 )]
            uint64_t   *pool;
    };
};
