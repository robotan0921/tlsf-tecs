
import("tTLSFStatistics.cdl");

[active]
  composite tTLSFMallocStatistics {
		
		entry sMalloc eMalloc;
		//call  siHandlerBody  ciBody;     /* 割込みサービスルーチン本体 */

		attr {
			ATR attribute = C_EXP("TA_STA"); 
			RELTIM cyclicTime = 4;
			RELTIM cyclicPhase = 1;
			size_t memoryPoolSize = 1024 * 1024;
		};

		cell tTLSFStatistics TLSFStatistics {
			cMalloc = TLSFMalloc.eMalloc;
			cMallocStatistics = TLSFMalloc.eMallocStatistics;
		};
		
		cell tCyclicHandler CyclicHandler {
			ciBody = TLSFStatistics.eiBody;
			attribute = composite.attribute;
	        cyclicTime = composite.cyclicTime;
	        cyclicPhase = composite.cyclicPhase;
		};

		cell tTLSFMalloc TLSFMalloc {
	    	memoryPoolSize = composite.memoryPoolSize;
	    };
		
		composite.eMalloc => TLSFStatistics.eMalloc;
	
	};