import_C( "t_stddef.h" );

signature sMallocStatistics {
	size_t getUsedSize(void);
	size_t getMaxSize(void);
};