/**
 *  VM1.cdl
 *
 */
import("EV3_common.cdl");

//[domain(HRP2, "trusted")]
//[domain(HRP2, "nontrusted")]
region rDomainEV3 {
	cell nMruby::tMrubyVM MrubyVM {

		mrubyFile = "$(MRUBY_LIB_DIR)/EV3_common.rb "
			"$(MRUBY_LIB_DIR)/RTOS.rb "
			"$(MRUBY_LIB_DIR)/Speaker.rb "
			"$(MRUBY_LIB_DIR)/Button.rb "
			"$(MRUBY_LIB_DIR)/Motor.rb "
			"$(MRUBY_LIB_DIR)/UltrasonicSensor.rb "
			"$(MRUBY_LIB_DIR)/GyroSensor.rb "
			"$(MRUBY_LIB_DIR)/ColorSensor.rb "
			"$(MRUBY_LIB_DIR)/TouchSensor.rb "
			"$(MRUBY_LIB_DIR)/LED.rb "
			"$(MRUBY_LIB_DIR)/LCD.rb "
			"$(MRUBY_LIB_DIR)/Battery.rb "
			"$(MRUBY_LIB_DIR)/Balancer.rb "
			"$(MRUBY_LIB_DIR)/SharedMemory.rb "
			"$(APP_RB)";
		cInit = VM_TECSInitializer.eInitialize;
		// cMalloc = TLSFMalloc1.eMalloc;
		cMalloc = TLSFStatistics.eMalloc;
	};

	cell nMruby::tMrubyTaskBody MrubyTaskBody {
      cMrubyVM = MrubyVM.eMrubyVM;
    };

	cell tTask MrubyTask1 {
	// 呼び口の結合
		cBody = MrubyTaskBody.eMrubyBody;
		//* 属性の設定
		taskAttribute 	= C_EXP("TA_ACT");
		priority 		= C_EXP("EV3_MRUBY_VM_PRIORITY");
		systemStackSize = C_EXP("STACK_SIZE");
		//userStackSize = C_EXP("STACK_SIZE");
	};

	cell tTLSFMalloc TLSFMalloc1 {
    	memoryPoolSize = 1024 * 1024;
    };
};

import("tTLSFStatistics.cdl");

region rDomainEV3 {
	cell tTLSFStatistics TLSFStatistics {
		cMalloc 		  = TLSFMalloc1.eMalloc;
		cMallocStatistics = TLSFMalloc1.eMallocStatistics;
	};

	cell tCyclicTask CyclicTask {
		cBody = TLSFStatistics.eBody;
        /*
		 *  TA_NULL     0x00U   デフォルト値
		 * 	TA_STA 		0x01U   周期ハンドラが動作している状態
		 */
		cyclicAttribute = C_EXP("TA_STA");
		cyclicTime 		= 4;
		cyclicPhase 	= 0;
		/*
		 * タスク例外処理ルーチンに指定できる属性はないため
		 * TA_NULLを指定する
		 */
		exceptionAttribute 	= C_EXP("TA_NULL");
		priority 			= C_EXP("EV3_MRUBY_VM_PRIORITY - 1");
		stackSize 			= C_EXP("STACK_SIZE");
	};
};
