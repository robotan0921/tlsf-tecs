import( <sMalloc.cdl> );
import( <sMallocStatistics.cdl> );

celltype tTLSFStatistics {
	require tKernel.eKernel;
	call 	sMalloc 			cMalloc;
	call 	sMallocStatistics 	cMallocStatistics;
	entry 	sTaskBody 		eBody;
	[inline]
		entry 	sMalloc 		eMalloc;

	attr {
		size_t 	maxSize = 1000000;
	};

	var {
		[size_is( maxSize )]int32_t *time;
		[size_is( maxSize )]int32_t *malloc;
		[size_is( maxSize )]int32_t *free;
        int32_t mallocNum;
        int32_t reallocNum;
        int32_t freeNum;
	};
};


/**
*	統計情報を取得するコンポーネントを加えた
*	TLSFコンポーネント
*/
[active]
composite tTLSFMallocStatistics {
	entry sMalloc eMalloc;

	attr {
		size_t 	memoryPoolSize 	= 1024 * 1024;
		/*
		 *  TA_NULL     0x00U   デフォルト値
		 * 	TA_STA 		0x01U   周期ハンドラが動作している状態
		 */
		ATR 	cyclicAttribute = C_EXP("TA_STA");
		RELTIM 	cyclicTime	 	= 1;
		RELTIM 	cyclicPhase 	= 1;
		PRI		priority		= C_EXP("EV3_MRUBY_VM_PRIORITY-1");
		SIZE	stackSize 		= C_EXP("STACK_SIZE");
	};

	cell tTLSFStatistics TLSFStatistics {
		cMalloc 		  = TLSFMalloc.eMalloc;
		cMallocStatistics = TLSFMalloc.eMallocStatistics;
	};

	cell tCyclicTask CyclicTask {
		cBody 			= TLSFStatistics.eBody;
		cyclicAttribute = composite.cyclicAttribute;
        cyclicTime 		= composite.cyclicTime;
        cyclicPhase 	= composite.cyclicPhase;
        priority 		= composite.priority;
		stackSize		= composite.stackSize;
	};

	cell tTLSFMalloc TLSFMalloc {
    	memoryPoolSize = composite.memoryPoolSize;
    };

	composite.eMalloc => TLSFStatistics.eMalloc;
};