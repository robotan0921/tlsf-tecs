
signature sMallocStatics {
	size_t getMaxSize(void);
	size_t getUsableSize(void);
	size_t getUsedSize(void);
	size_t getMallocSize(void);
	size_t getFreeSize(void);
	size_t getReallocSize(void);
};

celltype tTLSFStatics {
	require tKernel.eKernel;
	call 	sMallocStatics 	cMallocStatics;
	call 	sMalloc 		cMalloc;
	[inline]
		entry 	sMalloc eMalloc;
	[inline]
		entry 	siHandlerBody eiBody;

	attr {
		size_t 	maxSize = 1000000;
	};

	var {
		[size_is( maxSize )]
            int32_t *time;
		[size_is( maxSize )]
            int32_t *malloc;
		[size_is( maxSize )]
            int32_t *free;
        int32_t mallocNum;
        int32_t reallocNum;
        int32_t freeNum;
	};
};