import( <sMalloc.cdl> );
import( <sMallocStatics.cdl> );

celltype tTLSFStatics {
	require tKernel.eKernel;
	call 	sMallocStatics 	cMallocStatics;
	call 	sMalloc 		cMalloc;
	[inline]
		entry 	sMalloc eMalloc;
	[inline]
		entry 	siHandlerBody eiBody;

	attr {
		size_t 	maxSize = 1000000;
	};

	var {
		[size_is( maxSize )]
            int32_t *time;
		[size_is( maxSize )]
            int32_t *malloc;
		[size_is( maxSize )]
            int32_t *free;
        int32_t mallocNum;
        int32_t reallocNum;
        int32_t freeNum;
	};
};