/*
 *  tEV3Sample.cdl
 *
 *  VM$B$N8D?t$K1~$8$F(BCDL$B%U%!%$%k$rA*Br$9$k(B
 *  (VM$B$r#2$D;H$&>l9g!$(BVM2.cdl$B$r%$%s%]!<%H$9$k!K(B
 *
 */

import("VM1.cdl");
// import("VM2.cdl");
