import( <sMalloc.cdl> );
import( <sMallocStatistics.cdl> );
import( <kernel.cdl> );

celltype tTLSFMalloc {
    entry   sMalloc            eMalloc;
    entry   sMallocStatistics  eMallocStatistics;
    attr {
        /* memory pool size in bytes */
        size_t  memoryPoolSize;
    };
    var {
        [size_is( memoryPoolSize/ 8 )]
            uint64_t   *pool;
        size_t mallocSize;
        size_t freeSize;
        size_t reallocSize;
    };
};
