import( <sMalloc.cdl> );
import( <sMallocStatistics.cdl> );
import( <tCyclicTask.cdl> );

// const bool_t SEQUENTIAL = true;
// const bool_t TLSF_USE_SD = true;

celltype tTLSFStatistics {
	require tKernel.eKernel;
	call 	sMalloc 			cMalloc;
	call 	sMallocStatistics 	cMallocStatistics;
	call 	sDataqueue 			cDataqueue;
	[inline]
		entry 	sMalloc 		eMalloc;
	entry 	sTaskBody 			eBody;
};

celltype tSDTaskBody {
	call 	sDataqueue 	cDataqueue;
	entry 	sTaskBody 	eBody;

	attr {
		char *fileName;
	};

	var {
		// FILE *fp;
		int32_t *fp;
	};
};

/**
*	統計情報を取得するコンポーネントを加えた
*	TLSFコンポーネント
*/
[active]
composite tTLSFMallocStatistics {
	entry sMalloc eMalloc;

	attr {
		size_t 	memoryPoolSize 	= 1024 * 1024;
		char 	*fileName =	"/log.csv";
		uint_t 	queueSize = 1024;
		/*
		 *  TA_NULL     0x00U   デフォルト値
		 * 	TA_STA 		0x01U   周期ハンドラが動作している状態
		 */
		ATR 	cycleAttribute 	= C_EXP("TA_STA");
		RELTIM 	cycleTime	 	= 40000;
		RELTIM 	cyclePhase 		= 1000;
		PRI		priority 		= 9;
		size_t	stackSize 		= 4096;
	};

	cell tTLSFStatistics TLSFStatistics {
		cMalloc 		  = TLSFMalloc.eMalloc;
		cMallocStatistics = TLSFMalloc.eMallocStatistics;
		cDataqueue 		  = Dataqueue.eDataqueue;
	};

	cell tCyclicTask CyclicTask {
		cBody = TLSFStatistics.eBody;
        /*
		 *  TA_NULL     0x00U   デフォルト値
		 * 	TA_STA 		0x01U   周期ハンドラが動作している状態
		 */
		cycleAttribute 	= composite.cycleAttribute;
		cycleTime 		= composite.cycleTime;
		cyclePhase 		= composite.cyclePhase;
		priority 		= composite.priority;
		stackSize 		= composite.stackSize;
	};

	cell tDataqueue Dataqueue {
		dataCount = composite.queueSize;
	};

	cell tCyclicTask SDTask {
		cBody = SDTaskBody.eBody;
		/*
		 *  TA_NULL     0x00U   デフォルト値
		 * 	TA_STA 		0x01U   周期ハンドラが動作している状態
		 */
		cycleAttribute 	= C_EXP("TA_STA");
		cycleTime 		= 5000000;
		cyclePhase 		= 5000000;
		priority 		= composite.priority;
		stackSize 		= composite.stackSize;
	};

	cell tSDTaskBody SDTaskBody {
		cDataqueue = Dataqueue.eDataqueue;
		fileName = composite.fileName;
	};

	cell tTLSFMalloc TLSFMalloc {
    	memoryPoolSize = composite.memoryPoolSize;
    };

	composite.eMalloc => TLSFStatistics.eMalloc;
};