import( <sMalloc.cdl> );
import( <sMallocStatistics.cdl> );

celltype tTLSFStatistics {
	require tKernel.eKernel;
	call 	sMalloc 			cMalloc;
	call 	sMallocStatistics 	cMallocStatistics;
	[inline]
		entry 	sMalloc 		eMalloc;
	[inline]
		entry 	siHandlerBody 	eiBody;

	attr {
		size_t 	maxSize = 1000000;
	};

	var {
		[size_is( maxSize )]int32_t *time;
		[size_is( maxSize )]int32_t *malloc;
		[size_is( maxSize )]int32_t *free;
        int32_t mallocNum;
        int32_t reallocNum;
        int32_t freeNum;
	};
};


/**
*	統計情報を取得するコンポーネントを加えた
*	TLSFコンポーネント
*/
[active]
composite tTLSFMallocStatistics {
	entry sMalloc eMalloc;

	attr {
		ATR 	attribute 		= C_EXP("TA_STA");
		RELTIM 	cyclicTime	 	= 1;
		RELTIM 	cyclicPhase 	= 1;
		size_t 	memoryPoolSize 	= 1024 * 1024;
	};

	cell tTLSFStatistics TLSFStatistics {
		cMalloc 		  = TLSFMalloc.eMalloc;
		cMallocStatistics = TLSFMalloc.eMallocStatistics;
	};

	cell tCyclicHandler CyclicHandler {
		ciBody 		= TLSFStatistics.eiBody;
		attribute 	= composite.attribute;
        cyclicTime 	= composite.cyclicTime;
        cyclicPhase = composite.cyclicPhase;
	};

	cell tTLSFMalloc TLSFMalloc {
    	memoryPoolSize = composite.memoryPoolSize;
    };

	composite.eMalloc => TLSFStatistics.eMalloc;
};