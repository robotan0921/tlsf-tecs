/**
 *  VM1.cdl
 *
 */
import(<bridge.cdl>);
import("tTLSFStatistics.cdl");

cell nMruby::tMrubyVM MrubyVM {
	mrubyFile =
		"$(MRUBY_LIB_DIR)/RTOS.rb "
		"$(MRUBY_LIB_DIR)/LED.rb "
		"$(MRUBY_APP_DIR)/rtos_debug.rb";

	cInit = VM_TECSInitializer.eInitialize;
	cSerialPort = SerialPort1.eSerialPort;
	// cMalloc = TLSFMalloc1.eMalloc;
	cMalloc = TLSFMallocStatistics1.eMalloc;
};

cell nMruby::tMrubyTaskBody MrubyTaskBody {
   cMrubyVM = MrubyVM.eMrubyVM;
};

cell tTask MrubyTask1 {
// 呼び口の結合
	cTaskBody = MrubyTaskBody.eMrubyBody;
	//* 属性の設定
	attribute 	= C_EXP("TA_ACT");
	priority 	= 10;
	stackSize 	= 4096;
};

// cell tTLSFMalloc TLSFMalloc1 {
	// memoryPoolSize = 1024 * 1024;
// };
cell tTLSFMallocStatistics TLSFMallocStatistics1 {
 	memoryPoolSize = 1024 * 1024;
};